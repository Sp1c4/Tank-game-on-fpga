module DCU();

endmodule