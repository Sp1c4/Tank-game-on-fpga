module DCU_ctr();

endmodule